`define TLBP  3'b001
`define TLBR  3'b010
`define TLBWI 3'b011
`define TLBWR 3'b100
`define TLB_LINE 32
`define TLB_WIDTH 5
`define kseg0 3'b100
`define kseg1 3'b101
`define ASID 7:0
`define VPN2 31:13
`define ASID 7:0
`define GLOBAL 0
`define VALID 1
`define DIRTY 2
`define UNCACHE 5