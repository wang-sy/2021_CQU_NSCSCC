`include "defines.vh"

`define INIT_DECODE {8'b0, 3'b0, 1'b0, 5'b0, 1'b0, 5'b0, 1'b0, 5'b0}
`define ORI_DECODE {`EXE_ORI_OP, `EXE_RES_LOGIC, 1'b1, rt, 1'b1, rs, 1'b0, 5'b0}